`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Submodule Name: VGADisplayer
//////////////////////////////////////////////////////////////////////////////////

module VGADisplayer(
    //====================================================
    //=======           Input                       ======
    //====================================================
    input                   clk,        // 25 MHz clock
    input                   rst,        // Asynchronus reset
    input      [2:0]        car_state,  // RYG 1-bit encode  
                                        // Red/Yellow/Green light of car 1:on 0:off
    input      [3:0]        man_state,  // 1~8 Grenn light of man, 1-8: eight seperated motion, 
                                        // 0: red
    //====================================================
    //=======           Output                      ======
    //====================================================
    output reg [3:0] vgaRed,
    output reg [3:0] vgaBlue,
    output reg [3:0] vgaGreen,
    output     Hsync,
    output     Vsync
    );
    
    wire car_R, car_Y, car_G;
    wire [3:0] man_G_ID;
    wire man_R;

    assign  {car_R,car_Y,car_G} = car_state;
    assign  man_G_ID = man_state;
    assign  man_R = ~|man_state;


    //-----Value of light figure-------------------------
    //car black: R3-R0, G2-G0, B3-B0 all 0
    parameter [9999:0] black_G3       = 10000'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    //car red: B3-B0, G2-G0 all 0; R3-R0 the same
    parameter [9999:0] red_R3         = 10000'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter [9999:0] red_G3         = 10000'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    //car yellow: B3-B0 all 0; G3 all 1; R3-R0, G2-G0 the same
    parameter [9999:0] yellow_R3      = 10000'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    //car green: R3-R0, B3-B0 all 0; G3 all 1; G2-G0 the same;
    parameter [9999:0] green_G2       = 10000'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    //man redman
    parameter [22499:0] redman_R3     = 22500'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111001111111001111111001111111011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111001111111001111111001111111011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111001111111001111111001111111011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111001111111001111111001111111011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111001111111001111111001111111011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111001111111001111111001111111011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111001111111001111111001111111011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111000111111001111111001111111001111111001111111001111111011111110000000000000000000000000000000000000000000000000000000000000000000000000111111001111111000111111001111111001111111001111111001111111001111111011111110000000000000000000000000000000000000000000000000000000000000000000000000111111001111111000111111001111111001111111001111111001111111001111111011111110000000000000000000000000000000000000000000000000000000000000000000000000111111001111111000111111001111111001111111001111111001111111001111111011111110000000000000000000000000000000000000000000000000000000000000000000000000111111001111111000111111001111111001111111001111111001111111001111111011111110000000000000000000000000000000000000000000000000000000000000000000000000111111001111111000111111001111111001111111001111111001111111001111111011111110000000000000000000000000000000000000000000000000000000000000000000000000111111001111111000111111001111111001111111001111111001111111001111111011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111001111111001111110001111111001111111000000000001111110000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111001111111001111110001111111001111111000000000001111110000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111001111111001111110001111111001111111000000000001111110000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111001111111001111110001111111001111111000000000001111110000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111001111111001111110001111111001111111000000000001111110000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111001111111001111110001111111001111111000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111110001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111110001111111000000000001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111110001111111000000000001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111110001111111000000000001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111110001111111000000000001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111110001111111000000000001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111110001111111000000000001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter [22499:0] redman_R2     = 22500'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111001111111001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111001111111001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111001111111001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111001111111001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111001111111001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111001111111001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111001111111001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111001111111001111111000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111001111111001111111001111110011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111001111111001111111001111110011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111001111111001111111001111110011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111001111111001111111001111110011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111001111111001111111001111110011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111001111111001111111001111111001111110011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000111111001111111001111111001111111001111110001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000111111001111111001111111001111111001111110001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000111111001111111001111111001111111001111110001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000111111001111111001111111001111111001111110001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000111111001111111001111111001111111001111110001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000111111001111111001111111001111111001111110001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111001111111001111111001111111001111110001111111001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001000001000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111001111111001111111001111111001111111000000000001111110000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111001111111001111111001111111001111111000000000001111110000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111001111111001111111001111111001111111000000000001111110000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111001111111001111111001111111001111111000000000001111110000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111001111111001111111001111111001111111000000000001111110000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111001111111001111111001111111001111111000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111110001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111110001111111000000000001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111110001111111000000000001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111110001111111000000000001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111110001111111000000000001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111110001111111000000000001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111110001111111000000000001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111110001111111000000000001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter [22499:0] redman_R1     = 22500'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111110001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111110000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111110000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111001011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111001011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111001011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111001011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111001011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111001011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111001011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111001011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111001011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111001011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111001011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111001011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111001111111001111001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111001111111001111101001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100111110001111111001111111000111111001111110011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111101111101001111111001111111000111110001111111011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111001111111001111111001111111000111111011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111001111111001111111001011111001111111011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111001111111001111111001011111001111111011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111110001111111001111111001111111001111111011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000111101000111111001111110001111110001111111001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110001011111001111111001111111001111111001011111001111111001111111011111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111101001111111001111111001111110001111101001111111011111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111001111111001111111001011111001111111001111111011111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111001111111001111111001011111001111111001111111011111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111001111111001111111001011111001111111001111111011111110000000000000000000000000000000000000000000000000000000000000000000000001111111001101111001111101001111111001111111001111111001111111001111111011111110000000000000000000000000000000000000000000000000000000000000000000000001111111000011111000111110000111111001111111001111110001111111001111111011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111001111111000000000001111111001111111001111101000000000001111110001111100000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001011111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001011111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001011111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001011111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001011111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111110001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001011111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001011111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001011111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001011111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001011111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001011111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001111111000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000000111110000111111000000000001111111001111111001111111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111110001111111000000000001111111001111111001011111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001011111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001011111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111001011111000000000001111111001111110000000000000000000000000000000000000000000000000000000000000000000000001111110001111111000000000001111111001111111001111111000000000001111110001111110000000000000000000000000000000000000000000000000000000000000000000000000111110001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000111110001111111000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111001111111001111111000111111001111111000000000001111110000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111001111111001111111001111111001111111000000000001111110000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111001111111001111111001111111001111111000000000001111110000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111001111111001111111001111111001111111000000000001111110000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111000111111001111111001111111001111111000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000111110000000000001111111000111111001111111001111111001111111000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111001111111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001011111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001011111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001011111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001011111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001011111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001011111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111001111111000000000001111101000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111001111111000000000001011101001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001011111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001011111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001011111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111110001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001011111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001011111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001011111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001011111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001011111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001011111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111001111111000000000000111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000000000001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111101001111111000000000001011110001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110001111111000000000001111110001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111110001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111011111100001111111000000000001111110001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111011111110001111111000000000001011111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111011111110001111111000000000001011111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111011111110001111111000000000001011111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110011111100001111111000000000001011111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111010011100001111111000000000001011111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111110001111111000000000001011111001111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter [22499:0] redman_R0     = 22500'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000100000001010000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000100000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000100000001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001111111000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000111111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001001000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000011000000000000000001000000010001000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000100000010000000000000000000001000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100100000000000000010000001000100000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001000010001000000000000001000000001001000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100001001000000000000000000000001000100000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001100010000000000000000000000000001000000010000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000010000001000010000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000101100000000100001001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000001000010000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111001101111000000000000111111101111111000011101000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001001110001000000000001000000001111111001100001000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001000000000000000000111111000000000000111111000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000001000001001000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110001011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000111110001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001000000000000000000001000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000001000000100000000001100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100011000000000000000000000000010000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000001100001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001111111000000000001011111001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100011000000000000000000000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111011111110001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100010000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110011011110001111111000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    //man greenman1
    parameter [22499:0] greenman1_G3  = 22500'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111011111111100111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110011111011101111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111011111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110111111111111111111100000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110111111111111111111100000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111100000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110111111111111111111100000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110111111111111111111100000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110111111111111111111100000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111100000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110111111111111111111100000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110111111111111111111100000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111111111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111111111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111111111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111111111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111111111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111111111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111111111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111111111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111111111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111110000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000111111111011111111110000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000111111111011111111110000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000111111111011111111110000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000111111111011111111110000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000111111111011111111110000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000111111111011111111110000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000111111111011111111110000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000111111111011111111110000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter [22499:0] greenman1_G2  = 22500'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111100111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111101111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111101111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111011111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111110111111111000000000000010111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111101111111011111110100000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111100000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110111111111111111111100000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111100000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111100000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111100000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110111111111111111111100000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111101111111111111111111100000000000000000000111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111100000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000100100000110011111111100000000000000000000011111101000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000011111111101111111110000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000111111111111111111110000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000111111111111111111110000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000111111111111111111110000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000111111111111111111110000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000111111111111111111110000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000111111111111111111110000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000111111111111111111110000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000111111111111111111110000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000011111111011111111100000000000010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000111110110000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000011000111000001000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000010000011000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter [22499:0] greenman1_G1  = 22500'b000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011111111110011011101100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000011101000000010000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111100111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111110011111111110111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111111101111111110111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111110111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111111110111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111110111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001011111111111111111110111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000011101111111101111110001111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110011111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111011111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111111011111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110011111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111111111111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110111111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111110000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110011111111001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101101111110111111111000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111111011111111000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111111111111111000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111111011111111000000000010111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111111111111111000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111000000000010111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111101111111110011111111000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111111111111111100000000010111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101011111101111111101111111110100000000001001000010111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000001010000000100000001000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101111111110111111111100000000000000000001011111110100000000000000000000000000000000000000010000000000000000000000000000000000000000101111111110111111100111111110111111111100000000000000000000011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110111111101111111110011111111000000000000000000001011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111101111111110111111111000000000000000000001011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111101111111110111111111000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111100111111110011111111100000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111101111111110011111111100000000000000000001011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111101111111110111111111100000000000000000001011111111100000000000000000000000000000000000000000000000000000000000000000000001011111111011111111011111111010011111001111111110011111111100000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000100000000010000000000000000000000000010100000000010000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000011111111001111111110000000000011111111100000000000000000000000000000000000000000000000000000000000000000000001011111111100000000000000000000000000000011111111011111111110000000001011111110100000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000011111111011111111110000000000011111110100000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000011111111111111111110000000000011111110100000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000011111111011111111110000000000011111110100000000000000000000000000000000000000000000000000000000000000000000001011111111100000000000000000000000000000011111111011111111110000000001011111110100000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000011111111001111111100000000000011111110100000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000011111111111111111110000000000011111110100000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000111111110101110001100000000000101111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000010111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000010111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101111110000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000001100000000001000000110011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000001011111110100000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001111111111000000000000000000010000000000011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000001011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000111111110000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101111110000001001000000000000000000000000000000111110111011111101100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101000000000000000000000000000000000000000000000000111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000000000000000001000000000000000000000111111101000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000001000000000000000000000111111101000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000000000000000001000000000000000000000111111101000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000000000000000000011111111011111111101101111111000000000000000000000000000000000000000000000000000111000111110111110011000000000000000000000000000000000000000000000001011111111101111111110000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000001011111111111111111110000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000111111111101111111110000000000000000000000000000000000000000000000000000000000100000000011111111100000000000000000000000000000000000000000000000000000011111111101111111110000000000000000000000000000000000000000000000000000000000100000000011111111100000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000001011111111111111111110000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000111111111101111111100000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000101111100011111111110000000000000000000000000000000000000000000000000000000000000000000000000001110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter [22499:0] greenman1_G0  = 22500'b001111111011111111101111111111111111110101111111101111111100111111110111111111011111111111111111111111111100111111111001111111101111111110011111111100000000000000000000000000000000000000000101110111100011011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000101111111111111111110110000000000000000000000000010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111011111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000101111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000101111111110111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000101111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000101111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001111011000000000100000000100111111100111111111110111101110001111101000000000000000000011000000010000000000110001010000000000000100101000000000000000000000000000000000000000000000011111000111111100111111111100001111011100000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001011111110111111111100111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000111111111001111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001011111111111111111110111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001011111111111111111110111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001011111111011111111110111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001011111111111111111110111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111011101111111110111111111101111101000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100010000001111111111100111100000000001000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000101111111100111111110000000000000000000000000000010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001000000010111111111111011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001000110000111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000011111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000101111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000111111111111011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000101111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001000000000101111111110111111111000000010000000000000000000000000000000000000000100000000000000000000000000000000000000010000000000000000000000000000000000000000110011001000011111101100010110000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111110101110000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010111111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000100000000000111111110111111111100000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000100000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000010111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000010111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001000000000000000000110111111101111111111100000000000000000010000000000000000000100000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000111111111111111111111000000000100001000000000000000000000000000000000000000010000000000000000000010000000000000000000000000000000000000000000000000000001111101110000010100000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110111111111011111110111111111010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000110111111111111111110111111110111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111101111111111011111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110111111111011111111000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000010111111111111111111011111111111111111100000000001000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000010111111100111111110111111111111111111110000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000010111111101111111110111111111011111111110000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001000000000000000000010111111111111111110111111111111111111110000000000000000000100000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000111111110011111011101111111100000000011111111110000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000011111000111110010111111110000000000011110000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000111001011111101100000000010111111101000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000110111111111111111110111111111100000000001111111110000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000010111111110111111110111111111100000000010111111111000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000111111110111111110111111111100000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000111111111111111110111111111100000000010111111110000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000001000000111111100111111110011111111100000000000111111111000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000010011111111111111101111111111100000000000111111110000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000111011111111111111110111111111000000000000111111110100000000000000000000000000000000000000000000000010000001000000000000100000000001000000011101101111011000000000000000001000000001100000000011101000011011111110000000000010000000010000000000000000000010000000000000000000000000000000000000000010000001000111111100011111000111111101000000000000000000001101000000101000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110111111111111111111011111111000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110111111111111111111000000000000000000001011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110011111111111111111111111111100000000000000000000011111110000000000000000000000000000000000000000010000000000000000000000000000001000000010101111111110111111111111111111111111111100000000000000000000111111111100000000000000000000000000000000000000010000000000000000000000000000000000000000101111111111111111111111111111111111111100000000000000000001011111111100000000000000000000000000000000000000010000000000000000000000000000000000000000001111111110111111110111111111111111111000000000000000000001011111110000000000000000000000000000000000000000000000000000000000000000000000000000000100101111111111111111111111111111111111111000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111111111111111111111111011111111000000000000000000000111111110000000000000000000000000000000000000000010001001111011111001101111100000011111111111111111010111111000011111000000000001011111111011111110011100000000110110110011111111110111111110000000000000000000000000000000000000000001100001000110000000000000000001000000010100000000010000000010000000001110000010100000000000000000000000000000000000000000000000000000000000000000000001011111111000000000000000000000000000000011111111111111111100000000001011111110000000000000000000000000000000000000000010000000000000000000000000000000011111111000000000000000000000000000000011111111111111111100000000000011111111000000000000000000000000000000000000000010000000000000000000000000000001011111111000000000000000000000000000000011111111111111111100000000001011111111000000000000000000000000000000000000000010000000000000000000000000000001011111111000000000000000000000000000000011111111011111111100000000001011111111000000000000000000000000000000000000000010000000000000000000000000000001011111111000000000000000000000000000000011111111111111111100000000001011111111000000000000000000000000000000000000000010000000000000000000000000000000011111111000000000000000000000000000000011111111111111111100000000000011111111000000000000000000000000000000000000000010000000000000000000000000000001011111111100000000000000000000000000000011111111111111111110000000001011111111000000000000000000000000000000000000000010000000000000000000000000000001011111111000000000000000000000000000000011111111011111111100000000001011111111000000000000000000000000000000000000000010001111111011111111101111111011111111110111111111100111111101011110111100000001110001110010000110001101111101111111111011111111011111111110000101110110000000000000000000000000000000000000000000000000000000000000000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100011111111011111111101000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111111100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000011111111011111111100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000011111111011111111100000000001000000000100000000000000000000000000000000000000010001111111000000000101111111001011111110101111000010000000101000111111000000001111111111101011111110010011000111111111011111111110100000010000000000010000000000000000000000000000000000000000000000000000000000000000000000111111110000000000001110001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000010111111110000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000011111111100000000010111111111000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000011111111100000000010111111110000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000111111111000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000111111110000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000011111111100000000010111111110000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000111111110000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000111110000110000001100000000010010001001110001110000000000000000000000000000000000000000010000001111001001100100000000011000101000101000010100000010000111111100100000001100000000011000000111111111110011011110011110101110000000010000001000010000000000000000000000000000000000000000000000000000000000001000111111000000000000000000000000000001011111010000000000000000000000000000000000000000010000000000000000000000000000001000000000000000000000000000001111111110000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000111111110000000000000000000000000000001011111111000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001111111110000000000000000000010000000001011111111000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000001111111111000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001001111111111000000000000000000010000000011111111111000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000100000001001111111111000000000000000000000000000000011111111001000000010000000000000000000000000000010000000000000000000000000000000000000000000000000001000000001111111111000000000000000000000000000001011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000100010001000000000000000000000000000000001100001111011000011000000000000000000000000000000010000000000001001111110000000011100001010101011011000101111100000001001111010110000000000010111101111010110110111110101000000000110111100001000000000010000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000111111111000000000000000000000000000000010000000000000000000000000000001000000000000000000010111111100000000000000000000000000000000000000000000000000111111111100000000000000000000000000000010000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000001000000011111111100000000000000000000000000000010000000000000000000000000000000000000000000000000010111111110000000000000000000000000000000000000000000000100111111111100000000000000000000000000000010000000000000000000000000000000000000000100000000000111111110000000000000000000000000000000000000000000000000011111111110000000000000000000000000000010000000000000000000000000000000000000000100000000000111111110000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000001000111111110000000000000000000000000000000000000000000000000111111111000000000000000000000000000000010000000000000000000000000000001000000000100000010000111111110000000000000000000000000000000000000000000000000111111111100000000000000000000000000000010000000000000000000000000000001011000010101001100000000110001000000000000000000000000000000000000000000000000101111100101000000100000000000000000000010000001010001000111100000000101111111110101111111011101111100000000010010000001000000000010000000011000000010100111000101110111100100000010000001010010000000000000000000000000000000011111111111110011000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000010000000000000000000000000000000011111110111111111100000000000000000000000000000000000000000000000000000000000000000100011111111100000000000000000000010000000000000000000000000000001111111110111111111100000000001000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000001011111111111111111100000000000000000000000000000000000000000000000000000000000000000000001111111100100000000000000000010000000000000000000000000000011111111111011111111100000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000010000000000000000000000000000001111111110111111111110000000000000000000000000000000000000000000000000000000000000000010001111111100000000000000000000010000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000010000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000010000000000000000000000000000001100010101000000110010000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000000000010001111111001111111001000000001001111100111111111000011100101000001010010100010001111111110111111101000000000110000010111111110010000000010010000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000010000000000000000000000000000000000010000100000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000010000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001011101000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    //man greenman2
    parameter [22499:0] greenman2_G3  = 22500'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111011111111101111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111011111111111111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111011111011101111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111011111111100000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111111111111100000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000111111101011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111110000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000111111111011111111111111111110000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000111111111011111111111111111110000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000111111111011111111111111111110000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000111111111011111111111111111110000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000111111111011111111111111111110000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000111111111011111111111111111110000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000111111111011111111111111111110000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter [22499:0] greenman2_G2  = 22500'b000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110111111111100111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111101111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111011111111101111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111011111111100000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111101111111111111111100000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110111111111000000000000000000000001001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111011111111100000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110111111111100000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000001000100100100100001110011111111100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000000000001011111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000111111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000111111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000011110000100001100000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001110111110000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000100000000000111001011000000000000000000000000000000000000000000000000000000100110000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000111111111011111111111111111110000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter [22499:0] greenman2_G1  = 22500'b000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000011111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000110011111111110011111100100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001001001001101000000110000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111110111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111110111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111110111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111110111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111110111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111110111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111110111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111110111111100011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000000010000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110011111111011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111110011111111011111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110011111111011111111101111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111111111111111011111111100111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110111111111011111111100111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111011111111100111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111100111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111111111111111011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100111111110011111111001111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000100000000000000000000000000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110011111111000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110011111111000000000000000000001011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110111111111000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111111011111111000000000000000000001011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111111111111111000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111111011111111000000000000000000001011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110011111111000000000000000000001011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111111111111111100000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000111111101111111110100000000000000000000110110101011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110111111111100000000000000000000000000000101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110111111111000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110011111111000000000000000000000000000000101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110111111111000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110111111111000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111110011111111100000000000000000000000000000101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000111111100011111111000000000000000000000000000000011111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111110111111111100000000000000000000000000000101111111110000000000000000000000000000000000000000000000000000000000000000000000011111110110011011011011110001011111111011111111100000000000000000011011111110100000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000011111111001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000011111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000011111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000011111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000011111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000011111111001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111101010000000000000000001111111111101111111110000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111110000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110110000001100000000001000001110011111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000001011111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000001011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000001011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000011111111011111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000001111111001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110100000000000000000000000000000111100001011011110001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000100000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000010111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000110111011000000000000000000000000000000000000000000000110000110001110001000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000010111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000010111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000010111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001011111100000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000011111110011111111000111111101000110100000000000000000000000000000000000000000001111111101111011000000000000000000000000000000000000000000000000000001111111110111111111110011111100000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000111111110111111111110111111100000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000111111110111111111110111111110000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000111111110111111111110111111100000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000111111110111111111110111111100000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000111111110111111111110111111100000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000111111110111111111110111111100000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000001111111111011111111110111111100000000000000000000000000000000000000000000000000101111111110000000000000000000000000000000000000000000000000000000000000011111110011111111110111111100000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter [22499:0] greenman2_G0  = 22500'b011111111111111111111111111001111111110101101111101111111100111111110111111111011111111100111111111111111101101111111101111111110111111110111111111010100000000000000000000000000000000000000101111111110111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000111111111111111111011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000011111111111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000011111111111011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000111111111110111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000111111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000111111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110010100000000100000000110011111001111111111110111011111011111011010110000000100000001000000010000000000100000010000000000000000100010100000000100000000000000000000000000000001110110001110110110111011111000111111011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111101111111101111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000111111110111111111111111111101111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001111111111111111111110111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001111111111111111111110111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001111111111111111111110111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000111111111111111111110111111111111111111000000000000000000000000000000000000000000000000000000000001000000000000000000000100000000100000000000000000001111111111111111111110011111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000001000100000111011111111111010111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000100000000000000000000000000000111111111101111111110000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000001000000010111111111110011111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000111111111111111111111000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000011111111110011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000111111111110111111110000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000111111111111011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000111111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000111111111100111111110000000010000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000100110011010111111001110011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100011111100111111101110000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000100111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000100000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000001000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000001000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000110011111110111111111100000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111101111000000000100100000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111001011000010100000000010000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110011111111111111110101111111100111111100100000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000110111111101111111111111111111111111111101111111110100000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000111111111111111111011111111111111111110111111111100000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000111111111111111110111111111111111111111111111110000000100000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010011111111111111111011111111111111111111111111110001000001000010000000000000000000000000000000000000100000000000000000000000000000000000000000000000010111111100111111110111111111111111111111111111110111000000000101000000000000000000000000000000000000100000000000000000000000000000000000000000000000010111111101111111110111111111011111111101111111111000000000100110000000000000000000000000000000000000100000000000000000010000000001000000000000000000010111111111111111110111111111111111111101111111111000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111011011111000101111110100000000001100000000010010011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011001001100100111001110000000000000000000000100110000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110000011001101111101000000000000000000001111111100000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000110111111111111111111111111111100000000000000000000111111111000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010111111111111111111111111111100000000000000000001111111111000000100000000000000000000000000000000000100000000000000000000000000000000000000000001000010111111111111111110111111111100000000000000000010011111111000100000000100000000000000000000000000000100000000000000000000000000000000000000000000000010111111111111111110111111111100000000000000000001011111111010000000000100000000000000000000000000000100000000000000000000000000000000000000000000000000111111111111111110111111111100000000000000000000011111111000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111111111111101111111111100000000000000000000011111111010011000000000000000000000000000000000000100000000100000000000000000001000000000000000000010111111111111111110111111111000000000000000000001011111111010000001000000000000000000000100000000000100010000100000000110100000001100110000100001111010000000101000000001000000001100000000000000000000010110111101111111101001100000000000010100001001000000000000000000000000000000000000000000000000000000011111001001111000111111100000000000000000000000000000000010000000000000000000000000000000000000000000000000100000000000000000000000000000000000000010111111101111111111011111111000000000000000000000000000000001111111101000000000000000000100000000000100000000000000000000000000000000000000000000000010111111111111111111011111111100000000000000000000000000000101111111101000000000000000000000000000000100000000000000000000000000000000001000000000000010111111111111111111111111111100000000000000000000000000000001111111100000000000000000000000000000000100000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000101111111100000000000000000000000000000000100000000000000000000000000000000000000000000000010111111111111111111111111111100000000000000000000000000000101111111110000000000000000000000000000000100000000000000000000000000000000000000000000000110111111101111111101111111111000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111011111111100111111111100000000000000000000000000000111111111001000000000000000000000000000000000000000000000000000000000000000000000000001000000111111101111111111011111111000000000000100000000000000000001111111101000000000000000000000000000000110001010111110101111111000101100000001101111010111011011001011110000000000000001111111011000110011000000100001111110100001011110011010100100000000010000000000000000000000000000000000000000100000000000000000000000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000111111111100000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000111111111100000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000111111111110000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000111111111100000000000000000000011111111011111111110000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000111111111100000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000111111111100000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000111111111110000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000111111111100000000000000000000011111111011111111110000000000000000000000000000000000000000000000000000000000000111111011001111111111111110001111111110011111101010111111100011110111100000000100000000011000110001111111101101111111111111111100111111110100000111010000000000000000000000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000100100011111111001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111011111111110000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000011111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111111110000001001000000000100000000000000000000000000000000000000000111111110100000001111111110001111011110111111000000000000100000110111000000001111111111101110111111010001000101101111011111111110000000010100100000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000001000000001000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000011111111100000000000111111110000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000011111111100000000001111111110000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000011111111100000000000111111110000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000011111111100000000000111111111000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000011111111100000000000111111110000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000011111111100000000000111111110000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110100000000000111111110000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000110000100110000001100000000000100001001110011010001100011100000000000000000000000000000000100001110100001000111000000001100001100111100000100000000001111111111110000001100000000011100001111111111111101111111000011100110000000010101000100000100000000000000000000000000000000000000000000000000000000001000111111000000000000000000000000000001011111100101111111101000000000000000000000000000000100000000100000000000000000001000000000000000000000001000000111111110000000000000000000000000000000011111111001111111101000000000000000000100000000000100000000000000000000000000001000000000000000000000000000001111111110000000000000000000000000000000011111111101111111001000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000001011111111111111111101000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000001111111111011111111110000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000011111111111101111111100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000011111111101111111000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001111111101100000000000000000000000000001011111111001111111001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101000000000000000000000000000001110001100100000001111000001110000000000000000000000100000000100001111110100100101000011110101011000110101111000000000000011010110000000000000111101101011100001111011110011111111100011000011100000000000000000000000000000000000000000000000000000000000000000000000110110110100000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000001000000000000000000000000000000111111110100000000000000000000000000000000000000000000000011111111111000000000000000000000100000000000000000000000000000000000000000000000000000000000111111101000000000000000000000000000000011100000000000000011111111111000000000000000000000100000000000000000000000000000000000000000000000000000000001111111111100000000000000000000000000000100100000010000000011111111110000000000000000000000100000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000010111111110000000000000000000000100000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000100000000010111111111000000000000000000000100000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000111111110000000000000000000000100000000000000000000000000000000000000000000000000000000000111111110100000000000000000000000000000000000000000000000010111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111011100000000000000000000000000000000000000000000000010111111101000000000000000000000100000000100000111110000000001000111110011000000100001111001000000101000000001000000000000000000011000000001100000011011000010001011000010101001101100000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000011111111100000000000000000000000100000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000001111111111000000000000000000000100000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000010111111111000000000000000000000100000000000000000000000000001000000000000000000000000000000111111111000000000000000000000000000000000000000000000110000111111110000000000000000000000100000000000000000000000000001000000000000000000000000100001111111111000000000000000000000000000000000000000100000100011111111110000000000000000000000100000000000000000000000000001000000000000000000000000000000111111111100000000000000000000000000000000000000100000000000111111101000000000000000000000100000000000000000000000000001000000000100000000000000000001111111111000000000000000000000000000000000000000100000000011111111110000000000000000000000100000000000000000000000000000000000000000000000000001000000111111111100000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000111110010011111011000011000001100001000100000000000000000000000000000000000000001110010011110000001000000000000000000000111111111101111111111000000101011111111111111111010110011110000110100010100010001111111100111111111000000001111111111001111011000011100000110000000110000000000000000000000000000000111111111111111111110111111111000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000100000000000000000000000000001111111111111111111111111111111000000000000000000000000000000000000000000000000101111111100000000000000000000000000000000100000000000000000000000000001111111111111111111110111111101000000000000000000000000000000000000000000000000101111111100000000000000000000000000000000100000000000000000000000000001111111111111111111110111111111000000000000000000000000000000000000000000000000101111111100000000000000000000000000000000100000000000000000000000000001111111111111111111110111111011000000000000000000000000000000000000000000000000111111111110000000000000000000000000000000100000000000000000000000000001111111111111111111110111111111000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000100000000000000000000000000001111111111111111111110111111111000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000100000000100000000000000000000111111110011111111110111111110100000000000000000000000000000000000000000000000001111111100000000000000000000100000000000000000000000000000000000000001100110111100001000000011000011000000000000000000000000000000000000000000000000100011100101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    //man greenman3
    parameter [22499:0] greenman3_G3  = 22500'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111011111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111011111111000000000011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111011111111101111111000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000001111111111111111111011111111101111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000001111111111111111111011111111101111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000001111111111111111111011111111101111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000001111111111111111111011111111101111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000001111111111111111111011111111101111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000001111111111111111111011111111101111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000001111111111111111111011111111101111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000001111111111111111111011111111101111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000001111111111111111111011111111101111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000001111111111111111111011111111101111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000011111111101111111110111111101011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000011111111101111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000011111111101111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000011111111101111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000011111111101111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000011111111101111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000011111111101111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000011111111101111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000011111111101111111110111111111001111101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000001111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000001111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000001111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000001111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000001111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000001111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000001111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000001111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000001111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000001111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000001111111110111111111011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000001111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000001111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000001111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000001111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000001111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000001111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000001111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000001111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111011111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter [22499:0] greenman3_G2  = 22500'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110101111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111101111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111111111111110101111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101011111110011111111001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111101000000000001111111111101111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111110000000000000000000000101111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111101111111111111111100000000001101111111100111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000001111111110111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100111111111011111111100000000001111111111011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000111111111011111111101111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000001111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000001111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000001111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000001111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000001111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000001111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000001111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000001111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111101111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000111111100000111111011111111100011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000011111111111101111111100111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000011111111111111111111111111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000011111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000011111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000011111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000011111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000011111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000011111111111111111111011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000011111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001011111100000000000000000000000000000000111111100111111110011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000001111111110111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000001111111110111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000000000000000111111111011111111111111110110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110111111111000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110111111101000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111101111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter [22499:0] greenman3_G1  = 22500'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000001111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011111111110111111100100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111101111111110111111101101111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110001111111110111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111110111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111110111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111110111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111101111111110111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111110111111100111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110101111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100111111101111101011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110101111101101111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110111111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111110011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111101100000000111111111010111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111101000000000101111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110000000000001111111110111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110000000000001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110000000000001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110000000000001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111111000000000101111111100111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111100000000000011111111100111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111100001111101111111111011111111101011111111001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100111111110111111110100000000000011111101011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110011111111100000000000111111101111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111111111111111100000000000111111101111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111111011111111000000000010111111101011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111100000000010111111100011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111011111111100000000000111111101111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111111011111111100000000001111111101111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110111111111000000000010111111101111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110011111111000000000000111111100011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000000110000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000111111110011111111101111111101111111101011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000111111110011111111111111111111111111101011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000111111110111111111101111111110111111101111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000111111110111111111111111111110111111101111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000111111110011111111111111111111111111111011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000111111110111111111111111111111111111101011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000111111110011111111111111111111111111101111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000111111110011111111111111111110111111111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000001111111110011111111101111111110111111100011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101101111110011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111111111111110111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111110111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111110111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111110111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111111111111110111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111110011111110001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110111000000011111000000001111111001111111101011111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000101111111100111111101011111110111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000001111111111111111111111111111011111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000001111111111111111101011111110111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000001111111111111111101011111110111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000001111111111111111101011111110111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000001111111111111111101011111110111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000001111111111111111101111111111011111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000001111111110111111111111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000101111111100111111100011111110011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001010000000000000000000011111111101111111110000111111101111100100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000010111111101011111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000010111111111111111111111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000111111101011111110111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000001111111101111111110111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000111111111111111111111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000111111101111111111111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000111111100011111111111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000010111111110111111111111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000111111101011111110111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000001000000000100000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100111111110000000000000000000010111111100011111110111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110000000000000000000010111111101111111110111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111110000000000000000000000111111101011111110111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110000000000000000000000111111101011111110111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111111000000000000000000000111111101111111110111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111110000000000000000000000111111101111111110111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111110000000000000000000000111111101111111110111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110000000000000000000010111111101011111110111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111111000000000000000000001011111100010111110011111111010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111100111111110000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000000000000000000000000000001111111100111111100111111110000000000000000000000000000000000000000111111111010000000000000000000000000000000000000000000000000000000000000000000000001111111110111111100111111110000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000000000000000000000000000001111111110111111101111111110000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000000000000000000000000000001111111110111111101111111110000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000000000000000000000000000001111111110111111101111111111000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000000000000000000000000000001111111110111111100111111110000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000000000000000000000000000101111111110111111101111111111000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111100111111100000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001110111111000101111000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter [22499:0] greenman3_G0  = 22500'b000000000000000000000000000000000000000001111111100011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010111011111011100111011110011011110101001010101110111100111101110111111111001111111110111111101011111100111111111010111011100111101111011110010000000000000000000000000000000000000000000101110111100011010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111111111111111111000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111011110011110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000010000000100000001001011111101111111111110011001011011111101010110000000100100011000000000000000100110001110000000000000101001001001000000000000000000010000000000000000000111111111111111111101111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110101111111101111111101111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111011111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110111111111111111110000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110011111101101111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000100110000000001101111111010111100000000001000000000000000000010000000000000000000000000000000000000010000000000000000010000000000000010000000000000000000000000000101111111101011111110000000000000000000100000000010000000000000000000100000000000000000000000000001000000000000000000000000000000000000000000000000000001111111110011111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000101111111111111111111000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111110000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001111111100111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000010000000000010111111110100111100110000000101111110110001010100000000010100000111010010000100001011011000100110110000011000000000000000000000000000000000000000000000000000000000000000000000001000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110110101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000111111110111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000001011111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011111111111111111100000000000000000010000000000000000000100000000000000000000000000000000000000000000000010010000111100010000010000001011001000111110000000010000000011001101111111111111010000000101001000000100001101001110011110100100011010011111000000000000000000000000000000000000000000000000000000000111101011000000110000000110000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111111111111111011111110101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111101111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011111111111111111111111111001111111100000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111111111111111011111110111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111101111111111011111110111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111111111111110011111111101111111100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000010011111111111111111111111111111111111101000000000000000000100000000000000000000000000000000000000000000111111010011101000111110100110010010101001111110000000010100000011100000000000000000111100111000000000000111000101011111111110111010111011101000100000000000000000000000000000000000000000000000000000011011101000000000000000000110000000011000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111111111111110100000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111111111111111000000000101111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111111111111111000000000101111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000101111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111111111111111000000000101111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011111111111111111000000000101111111101111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111111111111101000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100011111100111111110110000000011001111100111111110100000000000000000000000000000000000000000000000000010000000000000000000000000001100001011010100000001100000001011001110111111111110110000010101111110000000000010000000010000000001000000010000000000000000000000000000000000000000000000000000000111111111001111101001111111000000000010001111111110101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011111101111111111111111111010000000010111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111110111111110011111110000000000010111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110111111111100000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110011111111000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111101111111110111111111010000000010111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011111111111111100111111110110000000010111111101011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111111011111111000000000000111111110011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000110011111111001111111010000000010001011110011111101100000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000110000100010000000000100000000100010010100000000000000000000000000000000000000000000000000000000000000000000000000000000101111111100000000000111111011101111111111111111011111111111111111011000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110000000001111111111011111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111011111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110000000000111111111111111111111111111011111111101111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110000000000111111111011111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111111111111111111111011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110000000001111111111111111111111111111111111111101111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000010000000001000000000111101111011111111100000000001000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000100011111111101111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011111111111111111101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111101000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011111111101111111100000100001000000000100000000000000000000000000000000000000000000011110010000011101111011000011111110111111110000000011101111110100010000000100000000001111111101011011000111111111011111111110100100001001000100000000000000000000000000000000000000000000000000000000000000001000000000001011110000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111110111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111100011111100100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000111000101100000001100000011101111111011101111000101111110011001001000000000000000000000000000000000000001110011001100000100000000000001000101001001100011010101000000011111000000110000000111100000000110101110111111111010111001110010000011000011000000000000000000000000000000000000000000000000000000000011111110000000000000000000001111111111101111110110101101111111101100000000000000000000000000000000000000000010000000000000000000000000000000000000010111111101000000000000000010101111111100111111100011111110011111111110000000000000000001000000000000000000000000000000000000000000000000000000000000010111111000000000000000000000101111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010111111110000000000000000000111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010111111110000000000000000000101111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000101111111110111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010011111110000000000000000000101111111110111111101011111110011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010111111110000000000000000000101111111111111111100011111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000011010100000000000000000000000000000011111111110111111110101111100100000000000000000000000000000000000000010010001110110000000000100101010100001111110100110111000000010011010010101111111010000000011100000000100000000011111001110110100001010000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000111111111100000101111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010111111110000000000000000000000000000000111111101111111110111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010111111110000000000000000000000000000010111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010111111110000000000000000000000000000010111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000010111111101111111110111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010111111100000000000000000000000000000010111111111111111110111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010111111100000000000000000000000000000010111111110111111110111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010011111110000000000000000000100000000001111111100111111110111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000011111001111111110000000000000000000010011010111111111101111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011100000000000000000000000001111001100111111110011110001010000000000000000000000000000000000000000000000000000000000000000000000000000000000111110101111110000000000000000000000000111111110011111111011111000100000000000000000000000000000000000000000000000000000000000000000000000000000000010111111110111111111110000000000000000001111111110011111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010111111101111111111000000000000000000010111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000010111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110100000000000000000011111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111111000000000000000000010111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010111111101111111111100000000000000000010111111111111111111111111111100000000000000000000000000000000000000000010000000000000000000000000000000000000010111111111111111111100000000100000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000110001110011111111011111110000000000000000000011100000011101000111110111101100000000000000000000000000000000000000000000000000000000000000000000000010000110000111111001000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111011111100010111010011110111100000000000000000010000000000000000000101111100110000000000000000000000000000000000000000000000000000000000000000000000101111111101111111111111111111100000000000000000010000000001000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000101111111110111111111111111111100000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000101111111110111111111111111111000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000101111111110111111111111111101000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000101111111110011111110111111110100000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000101111111110011111111111111111100000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110110000000000000000000000000000000000000011111111110000000000000000001000000000000000000000000000000000000000000000000000101111110000011111100011111101100000000000000000010000000000000000000110011011100000000000000000000000000000000000000000000000000000000000000000000000000000000000011111101000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111111111111101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011111110111111101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000011111111111111110100000000100000000010000000000000000000100000000000000000000000000000000000000000011110101001001011101011110010111111111101000110100111111110000101101010111111111111101101000011000111111010111111001011111111111100101110111101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    //man greenman4
    parameter [22499:0] greenman4_G3  = 22500'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000111111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000111111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000111111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000111111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000111111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000111111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000111111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000111111111111111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000111111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110100000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter [22499:0] greenman4_G2  = 22500'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111101111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111100111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111110111111111101111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111011111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111010000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111010111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000110011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111111111111110101111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110100000000000101111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001101111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001010000101011000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000010111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111011000000000000010111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter [22499:0] greenman4_G1  = 22500'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011111110101111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000101111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010001111111110111111111100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111110111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111101111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110111111111110111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111101111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000010000000011000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110111111111111011111101101111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000101110101111110001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110101111111101111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111100111111110011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000011111101011111001001111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000010001111111011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000111111101001111110111111111100000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000000100000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111101111110101011010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111110000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001111111110111111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110011111111001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000011111001101111110111111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111101000000000011111111011111111100111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101000000000011111111011111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101000000000011111111011111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101000000000011111111011111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000011111111011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000011111111001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101000000000011111111001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000011111111011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000011111111001111111100100111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000001000000000001010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000010111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000010111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110101111010100101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101111100000000001110111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000010111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110100000000010111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000010111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000010111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000010111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000100100000000001101000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter [22499:0] greenman4_G0  = 22500'b000000000000000000000000000000000000000000010010000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010111011111111111111011110011011010100101111101010111111101101101111101011001111111110111111111011101100101101111001011011100111101110111111010100000000000000000000000000000000000000000101110111100101010000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000000000000000000000000000101111111110111111110110000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000001111111110111111100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000001000000000000000000101111111110011111111000000000000000000000000000000000000001000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000101111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110011111110000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010001111000010000000100000000110101111101111111111111011011110001011111000000001000000000011011000010000000000100000010000000000000100000000100000000110000000000000000000000000000000011111111111111111101111111111101111111100000000000000000010000000000000000000100000000000000000000000000000000000000010000000000000000000000000000000111111111101111111100111111101111111111000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000011111111101111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110011111111111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110111111111111111111010000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000011111111101111111110111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000111111111111111111110011111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000011111111111111111110111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100011111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000000000000000100110000001001111111101110111100000000000000000000000000000000000000000000000000100000000000000000010000000000000000000000000000000000000000000000000000000000000101111111101001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000101111111110011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000111111111110111111110100010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000111111111110011111111000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000011111111110111111110000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000101111111100111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000101111111110011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000001111111100111111111100000010000000000000000000000000000000000000000000000000000000000000000000000000000000010000110000010000001011000000000111111111110000101101010000011101110111110001010000000000010110000111010000000110000111011100000110110001011100100000010000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111010110110110000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000110001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000100000000001111111110111111111100000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000001000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000100000000000000000000000000000000000000010000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000011111111101111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011111100111111111000000000000000000000000000000000000000100000000000000000000000000000000000000010000100010010010111101010000010000001000001001111111100000011010000001001111110000000000010001001111011000000100000001001110011110110000010101011111110000000000000000000000000000000000000000000000000001000111100010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100011111011111111110100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000011111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111111111111111011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001111111111111111110011111111100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000011111111100111111110111111111100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000011111111111111111110011111111100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000001000000000000000000000000000011111111111111111111111111111100000000000000000000000000000100000000000000000000000000000000000000010000110111010011101101110010100110100010101011011111100000000100000110010000000111111111110111111111011111100111110101011111111110100111110111111100100000000000000000000000000000000000000000000000000000011011100001111010111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000011111111111101111101111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011111111111111110111111111100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000011111111111111111110111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111111111111110111111111100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000011111111111111111110011111111100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000011011111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000011111111111111111111111111111100000000010000000000000000000100000000000000000000000000000000000000010000000000010000000001000000000010000001100000101000000000011010000001000000001000000000010000000001000000000100001000000000000010101000000100000000010000000000000000000000000000000000000000000000000001000000001011111010111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001111111111011111111000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001111111110011111111110000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000001111111110111111111100000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000100000000000000000000111111110111111110100000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000001000000001111111101111111111110000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001001111101001111111110010000000000000000000000000000000000000000000000000000000000000000010001001000011110101101111100010111100011101100000100110010111000000010100000000001111111011111000011000000010110101101011101111110111000110110110000000000000000000000000000000000000000000000000000000000000000001000000000101000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001111111111011111111101111111100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000001111111111011111111101111111100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000001111111111111111111111111111100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000001111111111011111111101111111100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000001111111111111111111101111111100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001101110101111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111001111110101111111110011011111011111111101100111101000000001110000000010100101110010100001111111100101110110001111011110101111100110101111110000000000000000000000000000000000000000000000000000000000001001111011111111111111111111100000000000000000000000000000000000000000000000000000000000010000000000010000000000000000000000000000000000000001000000001111111110111111111001111111101001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110011111111111111111100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000001111111110011111111111111111100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000001111111111111111111111111111100000000000000000000000000000000000000000000000000100000000010000000000000000000000000000000000000000000000000000000000001111111110011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001111111110111111111011111111110000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000010000000001100101111111110111111111100001110110000000000000000000000000000000000000000000000000010000111010010000011101111011000011001100111110010111111111010001111000010000000100000000001100110111011111000101100110011111111110100000010101000100010000000000000000000000000000000000000000000000000010111111010000000000011111111101111111111001010000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001111111110100000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000011111111111111111111111111110000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000011011111110000000000011111111111111111011111111110000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000011111111111000000000111111111111111111111111111111000100000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000011111111111000000000011111111111111111111111111110000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000011111111110100000000111111111111111111110111111110100000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000011011111101000000000011111111111111111111111111101000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001111111001000000000011101010101111111111010111101000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000000100011101000000000011010100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000010001111010000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000000000000000000011111111100000000000111111110000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001001000000000100000000011111111100000000010111111111000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000111111111100000000010111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111110000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000011111111100000000010111111110000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000011111110100000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000011111111100000000000111111100000000000100000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000111111110000001001010111111110000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000100000000010000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000111111111011111111111111111110000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000000011111111011111111111111111110000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000000111111111111111111110111111110000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000010010111111111111111111111111111110000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000000011111110111111111111111111110000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000000011111111111111111111111111110000000000100000000000000000000000000000000000000010000001010010010111101000000010000111111000000000001000000101000000100101110101111010100111000000001100000000100001111001100001110110100010101001000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110001101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000100000000000000000000000011111111101000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000000000000100000000000010111111100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000000000000000000000000010111111110000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000000010000000000000000000111111110000000000100000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000010010000000000000000001111111100000000000100000000000000000000000000000000000000010000100110011011111101100011000111110010101100010111111101101110000010101100110011111111101001000001100000000111001001011110111110000100110111010100110000000000000000000000000000000000000000000000000000000000000000000000011111110100000000001111111101000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000100011111111010000000001111111100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000000111111111110000000001111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000010111111111110000000001111111110110000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000111111111100000000011111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000010111111111000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000111111110000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000000011111111110000000010111111110000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000010111111100000000011000001010100000000000000000000000000000000000000000000000010000000000010000000001000000000010010101000000000001000000001000000010111010100100000000011100000101001000100100001000000000000010100000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000010000000000010000000000000000000000000000000000000001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000000000000000000000000000000000000001000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000001000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000010000000000010000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    //man greenman5
    parameter [22499:0] greenman5_G3  = 22500'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111011111111101111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111101111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111011111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111011111011101111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111011111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111011111011111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111011111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111011111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111011111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111011111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111011111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111011111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111011111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111011111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111011111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111110000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000111111111011111111110000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000111111111011111111110000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000111111111011111111110000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000111111111011111111110000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000111111111011111111110000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000111111111011111111110000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000111111111011111111110000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000111111111011111111110000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter [22499:0] greenman5_G2  = 22500'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111100111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111101111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111011111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111101111111111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111011111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110111111111011111110100000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111101111111111111110100000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111100000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111100000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111100000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111100000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111100000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111100000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111100000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000100100000110011111111000000000000000000000011111101000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000011111111101111111110000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000111111111111111111110000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000111111111111111111110000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000111111111111111111110000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000111111111111111111110000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000111111111111111111110000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000111111111111111111110000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000111111111111111111110000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000111111111111111111110000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000011111111011111111100000000000010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001111110110000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000011000111000001000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000010000011000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010;
    parameter [22499:0] greenman5_G1  = 22500'b000000000000000000000000000000000000000011111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000011101000000010000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111100111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110011111111110111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111110111111101111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111110111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111001111111110111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111001111111110111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101111111101111110011111110011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001000001010000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000111111011111101111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111110011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111110111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111011111111110000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110011111111101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110111111111000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110111111111100000000000111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111111111111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111111111111111000000000000111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111111011111111100000000000111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111100000000010111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111111111111111100000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111111111111111100000000010111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110011111111100000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000001000000000100000001000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110101111110111111110111111110100000000000000000000111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110111111100111111110011111111100000000000000000000011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111100111111110011111111100000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110111111100111111110011111111100000000000000000001011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110111111100111111110111111111100000000000000000001011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111100111111110011111111100000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111100111111110011111111100000000000000000000011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111101111111110111111111100000000000000000001011111111100000000000000000000000000000000000000000000000000000000000000000000000011111111011111111011111111011011111001101111110111111111100000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000100000000010000000000000000000000000010100000000110000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000011111111101111111100000000000011111110100000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000011111111111111111110000000001011111110100000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000011111111101111111100000000000011111110100000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000011111111111111111110000000000011111110100000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000011111111111111111100000000000011111110100000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000011111111101111111110000000001011111110100000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000011111111101111111100000000000011111110100000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000011111111111111111110000000000011111110100000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000111111110001011101100000000000101111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000010111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101111110000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000001000000000001000001110011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000001011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000001011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000001011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000001011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000111111110000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101111110000001001000000000000000000000000000000111110111011111101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000011111111010000000000000000000000000000000000000000000000000000000000000011111111011111111101101111110000000000000000000000000000000000000000000000000000111000111110111110010000000000000000000000000000000000000000000000000011111111101111111110000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000011111111101111111110000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000011111111101111111110000000000000000000000000000000000000000000000000000000000100000000011111111100000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000111111111101111111100000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000101111100011111111110000000000000000000000000000000000000000000000000000000000000000100000000001110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000001000;
    parameter [22499:0] greenman5_G0  = 22500'b001101111011011111100111111110011111110101111111101111111110101111110111111011011111111110001111101011111100111111111001111111101111111111000101111100000000000000000000000000000000000000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000101111111111111111111100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111111011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111011111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110111111101100000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000111111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000111111100111111111100011111011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110111111111100111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111001111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111011111110111111110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110111111111111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111011111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000011111010101111111110111111110111111101000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100010000001111111111110111100100000001000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000011000000001110111111100111001100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111111111011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111111000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111011111111000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111001000011111101110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010000000010000000000010111111110000111110000000000101111100100000110100000000010000000111000100010110001011011001100110100000001001010010000000000000000000000000000000000000000000000000000000011110111111010101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111101111111111000000000100000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000100000100000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111101111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111111111111111000000000100001000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000111101110000010100000000110000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110111111111011111110111111111011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111111111111100011111111111111111101001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111101111111111011111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111101111111111011111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111111111111111011111111111111111100000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111101111111110111111111011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111111111111110111111111111111111110000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110011011011101111111100000000011011011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111001111110010111111110000000000011110000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110001011001011111101100000000010111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111111111111101011111111000000000010111111110100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111111111111110111111111000000000010111111101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110111111111100000000010111111110100000000100000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000111111111111111110111111111000000000010111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000111111101111111110111111111000000000000111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111110111111110011111111100000000010111111101000000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000111011111111111111110111111111000000000000111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001110011111111011111001111111000000000000010010010001110100010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001000111111101001111000111111111100000000000000000001101000000101000000000000000000000000000000000000000000000000000000000000000000000000000000011111101100001111101001111111011111110010000000000000000001111100110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111000000000000000000001011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110111111111111111111111111111000000000010000000001011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110011111111111111111111111111010000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111111111111011111111000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111111111111111111111000000000000000000001011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110111111111111111111111111110000000000010000000001011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111111111111110111111111011111111000000000010000000000111111110010000000000000000000000000000000000000000001101010010111101101110100001011111111111111111010111111001011111000010000001001111111011111000001100000000110110101011011111110110111111000000000000000000000000000000000000000000100001000110000000000000000000000000010100000000010000000010000000001110000010100000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000011101111111100011110000000001011111111000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000011111111111111111100000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000011111111111111111110000000001011111111000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000011111111111111111100000000001011111111000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000011111111111111111110000000001011111111000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000011111111111111111100000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000011111111111111111110000000001011111111000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000011111111111111111100000000001011111111000000000000000000000000000000000000000000001111111001111111100111111010111111110111111111100101111100011110111100000001110100010010000111001101111101111111111011111111111111111111000101110100000000000000000000000000000000000000000000000000000000000000000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111101000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111100000000001000000000100000000000000000000000000000000000000000000111011011000000101111111000011011110101111000010000000100000110111000000001111111111101011111100011011000111010111011111111110100000011000000000000000000000000000000000000000000000000000000000000000000000000000000000101011110000000000001110000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000010111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000010111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000010111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000010111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000010111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000111111100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000111110000111000001100000000010010000001110001110000000000000000000000000000000000000000000000001110011001100100000000010000101000101100010100000010001111111100100000001100000000011000001111111111110011001110011010101110000010011010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001111111110000000000000000000000000000000011111111000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111111110100000000000000000010100000000011111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000010000000001011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000010000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000111111111000000000000000000010000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001000111111111000000000000000000000000000000011111111001010000010000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001111111111000000000000000000000000000001011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000101000001000000000000000000000000000000001100001111011010011000000000000000000000000000000000000000000011001110110001000010100001010101011011000101111100000001001111010110100000000010111100101010110110111110101000100001110110100001000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000100010000010000000000000000000000000000000000000000000000000000000000000000000000000000000010111111100000000000000000000100000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101000000000000000000000000000000000000001011000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010111111110000001000000000000000000000000000000000000000100111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000100000000111111111100110000000000000000000000000000000000000000000000000000000000000000000100000000000111111110000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000001000000000101000111111110000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000100000010000111111110000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000011000010101101100000000110000000000000000000000000000000000000000000000000000101111100101000000100000000000000000000000000001010011000111100000010100111111110101111111011101111101001000010010000001100000000010000000001010000010100111000101110111100101000011010001010000000000000000000000000000000000011111111111110011000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000011111110111111111100000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000011111111111111111100000000001000000000000000000000000000000000000000000000000100000000011111111100000000000000000000000000000000000000000000000000000011111111111111111100000000001000000000000000000000000000000000000000000000000000000100001111111100100000000000000000000000000000000000000000000000010111111111011111111100000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000111111110111111111110000000000000000000000000000000000000000000000000000000000000000010001111111100000000000000000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000100000000011111111100000000000000000000000000000000000000000000000000000100010101000000110010000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000000000101111011111111001000000000001111100111111111000011100100110001010010100010101111111110111111101010110000111001110111111110010000000011000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001111101000000000000000000000000000001000010000000100000000010000100101100000010100100010000000000010000000000000000000010000000001010000000110000110010000000001100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000100000000010000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000011100011001000110100111010010111101111001101000110101000001100001010111111111111111111101000000000011101010011110001001110111111100001010111010100100;
    //man greenman6
    parameter [22499:0] greenman6_G3  = 22500'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter [22499:0] greenman6_G2  = 22500'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111111101111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111111100111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111111111111111101111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111100111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100011111110011111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111101000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000101111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100011111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101100000000000000000000001011101000100000000100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter [22499:0] greenman6_G1  = 22500'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010011111111111011111101100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111110111111110101111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111101111111100111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111001111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111001111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111101111011111111110000111101011101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000111110111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110101111101011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100111111110011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111111001111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000111111111000111111100000010001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100111111101000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100111111110000000000101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100111111110000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100111111101000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100111111100000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111100000000001011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111011111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000011111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111101001111110000000000001011101110000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000110000000100000000000000000001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111100000000000111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111100000000000111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111100000000000111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111100000000000111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111100000000000111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111100000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111101101111111101111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110011111110001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000011100000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111100000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101000000000000000000101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111100000000000000000000101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111010010000000000000000000010100010100011111110001111100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111101111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100111111110000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100111111111000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110000000000000000000000000000001000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111111000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001011111100111111111000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111101111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000100000000000000000000000000000110111110100111101000000000000000000000000000000100000000000000000000000000000000000000100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter [22499:0] greenman6_G0  = 22500'b000000000000000000000000000000000000000000010001000001101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001110111100011010101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111110011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111110011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111110111111101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000010100000100000000111001111101101111111110001001100011111101010100000000000000011100000000000000100110000110000000001000001000001010000001000010000000010000000000000000000011111111011111111101111111100111111111100000000000000000010000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000111111110111111111101111111100111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000011111111111111111110011111101111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000011111111111111111110111111111111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000011111111001111111110111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000111111111111111111110011111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000011111010001111111111011111111111111111100000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111110011111101001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000100110010000101101111110011111110100010000000000000000000000010000000000000000000100000000000000000000000000000000000000000010000000010000000000000000000000000000001111111101101111110000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000001111111100111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000010000011111111110111111111100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111110111111110000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111110011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111111111111110100000000000000000100000000000000000000000000000100000000000000000000000000000000000000000010000000010000000011010000000010011111010000111111111000000111111111110000010100000000010000000111010110010110001010001011100100110000111000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000111111111111111111111000000000100000000000000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001011111110111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001111111111111111111000000000100000000000000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001011111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011111111100111111101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111111101111011000000000000000000000000000000000000000000000000000000000000000000000000000000010001100011010111101001000010000000011000001111111000000011000000011101111111000000000010010001101001000000000001111001100011100101000101000011111000000000000000000000000000000000000000000000000000000011111110011111111011111110000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001111111111111111111011111111000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010111111111111111111111111110100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011011111111111111111011111111000000000010000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001111111111111111111011111111000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011111111101111111111011111111000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011011111110111111110011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110010111100010100010100011100010000000000000000000000000000000000000000000000000000000000000010101011010001011001110111110110111010010001011110000000010110000001100000000111111111011110000001111111000111111100001111111100111000101101111001000000000000000000000000000000000000000000000000000000011000110011111111100000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011111111111111111111000000000101111111100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011111111111111111111000000000101111111100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001111111111111111111000000000101111111100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011011111110111111111000000000101111111100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011111111111111111111000000000101111111110000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000000000011111111110111111110000000010101111111101000000000000000000100000000000000000000000000001000000000000000000000000000000000000000000000000000000000000001101111001011111100111111110111111111000100010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000011100100000000000000000011100000001000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001111111101111111110000000000011011111111000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000001111111110111111111010000000010111111110000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000000111111110011111111000000000010111111110000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000001111111110111111111100000000010111111111000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000000111111110011111111000000000010111111110000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000111111110011111111000000000010111111100000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000111111100011111110000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000011111110111111111000000000000111111110000000000000000000000000000000000000000000000000000011001101010111111101111101010111101010000000000011010000111000000011100000001111111111001110010011000000100111110100011011111100110101101100010000000000000000000000000000000000000000000000000000000000000000001000001000110000100100000000001000000101000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000001111111111111111111000000000010111111110000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000001111111111011111111000000000010111111110000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000001111111111111111111000000000010111111100000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000001111111111111111111000000000010111111110000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000001111111111011111111000000000010111111110000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000001111111111011111111000000000010111111110000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000001111111111011111111000000000010111111111000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000001111111111111111111000000000010111111100000000000000000000000000000000000000000000000000000011111110001011111101111111100011111111001111111101101111101111111110100000110011111111011111111110111100000111111111001111110101110111101100101111100000000000000000000000000000000000000000000000000000000000000000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000000000000000100011111111111111111100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111101000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000000000000000011111111111111111101000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000000000000000011111111111111111100000000000000000000000000000000000000000000000001000000000000010000000000000000000000000000000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000001111111101111111100000000000000000000000000000000000000000000000000000000000000010111111010000100101111101000001011110011111000011000011100111111100000000000100000000000000101001011110000111010110011111111100000001101000000000000000000000000000000000000000000000000000000000000000000000001001111111111111111001111111110000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001001000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000001111111111011111111111111111100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001111111111011111111111111111100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000001111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000001111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000101110011101001110011101111111000000000000000000000000000000000000000000000000000000000000000010000111011000100101000000000010000000001000001100111111111000010011100000000110000000110000000001000000000110000110001000001100000000101010001000000010000000000000000000000000000000000000000000000000110111110000000000000000000101111111100000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000000000011111111101000000000000000000111111111101000000001000000000100000000000000000000000000001000000000000010000000000000000000000000000000000000000000000011111111101000000000000000000101111111100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011111111110000000000000000000111111111101000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011111111110000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001111111110000000000000000000101111111101000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001111111111000000000000000000101111111111000100000010000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011111111110000000000000000000011111111110010000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111010000000000000000000001011011000111101000001001110000000000000000000000000000000000000000000010000001011000110111010010000110111110000000011000111010001111111010000110110100100010111011111101001111101000000010000010101100110110111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100111111111100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000010000000000000000000000000000000000000000000010001000000000000000000000000000000000000011111111101111111111000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111111000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000000000000000000000000000000000010111111110111111111000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111110111111111101100000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000010000000000100000000000111111101111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101100110110010000000000000000000011000100011000000010110011101000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000100010000000000000000000010000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101111101111111000100000000000000000000000000000000000000101110110010000000000000000000000000000000010000000000000000000000000000000000000000000000011111111111111111110110000000000000000000000000000000000000111111111100000000000000000000000000000000010000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000100000000000000011111111100000000000000000000000000000000010000000000000000000000000000000000000000000000011111111110111111111100000000000000000000000000000000000000011111111000000000000000000000000000000000010000000000000000000000000000000000000000000000001111111110111111110000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000011111111100000000000000000000000000000000010000000000000000000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000011111111100000000000000000000000000000000010000000000000000000000000000000000000000000000011111111101111111110100000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001011111110000000000000000000000000000000000000000111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010011100000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000100000101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000111111111100000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001111111111100000000000000000000000000000000000000111111111100000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000111111111100000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001111111111100000000000000000000000000000000000000111111111100000000000000000000000000000000010000000000000000000000000000000000000000000000000000100001111111110100000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111100000000000000000000000000000000000000111111111110000000000000000000000000000000000000000010000000000000000000000000000000000000000000000100111111010100000000000000000000000000000000000000011111111000000000000000000001000000000000000000000000000000000000000000000000000000000000000001111101011111001000000000000000000000000000000000000000101111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000001000000000000000000000000000001111111111111111111000000000000000000000000000001000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011111111111111111110010000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011011111110111111101110000000000000000000000000000000000000000000000000000000000000000000000000100000010000000000000000000000000000000000000000000000001011111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000000000001011111111111111110100000000100000000010000000000000000000100000000000000000000000000000000000000000001111001001100100101011010010111111111011001010000111111110000111111111110111101111111101100100001011100010111110001001110111101100001100010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    //man greenman7
    parameter [22499:0] greenman7_G3  = 22500'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111011001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter [22499:0] greenman7_G2  = 22500'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111111111111111101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111110011111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110100000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111100000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110100000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110100000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010001000111111110011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111100000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter [22499:0] greenman7_G1  = 22500'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100001010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010011111111111111011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111001111111110111111111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110111111111111111111111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111001111111110111111111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111001111111111111111111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111001111111111111111111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111111111111111111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111001111111111111111111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010011000000010000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000111110001111110101111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111111111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111110011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000111111111000111101000000010101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111110100000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110100000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110100011111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110101111101101111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110110111111111101111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111101101111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111111101111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111110111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111100111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000110000000000000000000001101001111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001000000000000000000000000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010111111110111111111000000000011000011100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110100000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110100000000000000000000111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110100000000000000000000111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110100000000000000000010111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111100000000000000000010111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110100000000000000000000111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110100000000000000000010111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100111111111000000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110100000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110100000000000000000000111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110100000000000000000010111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000010111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110100000000000000000000111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110100000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110100000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000010111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000001011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000010111111100111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter [22499:0] greenman7_G0  = 22500'b000000000000000000000000000000000000000001110001000011101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000111111100011010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111110011111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111011111101110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000010000000000000111001111101101111111110011101110001111111110100000000100010011010000000000000100101000110000000001000101001100000000010100010000000000000000000000000000011111111111111111100111111111101111111000000000000000000010000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000011111111001111111110111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000111111111111111111110111111111111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000111111111111111111110111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000111111111101111111110111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000011111111111111111110011111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000111111010001111111110011111111101111111000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111101010111111100011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000011011111000010111011100000110000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111101111111110000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000001111111110011111111000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111110011111111000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111110111111110000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111110011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000011111101100010110000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000111000000100010111111010000111101010000001101111111010000110000000000010000000111010000000110001010011101000110110100011000000000000000000000000000000000000000000000000000000000000000011111111111111110110000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000110011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001011111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001111111100111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001011111111111111111000000000000000000000000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001011111111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110111111111111011010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010011101111000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111110011111111011111111100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001111111111111111111111111110100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010111111111111111111011111110100000000000000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011011111111111111111011111111100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111111111111110100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000001000000000000000000000000000011111111111011111111111111111100000000000000000001000000000100000000000000000000000000000000000000000010001010010100110101110011110110011010001101011111000000000110000011100000000011111111011110000001011001000111001111011111111110111001010001101000100000000000000000000000000000000000000000000000000000011111100010000000000000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000110011111111100000000001111111111000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011111111111111111111000000000011111111110000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011111111110111111111000000000001111111110000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011111111111111111111000000000001111111101000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011111111111111111111000000000001111111101000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011011111111111111111000000000001111111101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011111111111111111100000000001111111100000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000000000011101111111111111110000000010001111111100100000000000000000100000000000000000000000000000000000000000010000000010000000001000000000000001000000001100001011110111000000001101111111111111111110111000101000000000100000000000000000110100000000000000010000000000000000000000000000000000000000000000000000000000000001110011110100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000000000000000000001111111110011111111010000000000000000001000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000111111110111111111010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000001111111110111111111100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000110111111110011111111100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000110000000100001111111110011111110100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000111111100011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000110101111101001111101100000000000000000000000000000000000000000000000000000000000000000000000011101101011100101101111101010111111010000000011111001011101000000011000000001111111111111000110101011111010110100101010110011110111111110000000000100000000000000000000000000000000000000000000000000000000000000100001000010000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000000000010111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111111100000000000000000000000000000000000000000000000000000000000000000000000011111111001001110101101111110011111111001111011100101110111000000000010000000010101111110111111101001111100101111111011111111111110111110000011110100010000000000000000000000000000000000000000000000000000000001001111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000000011111111111011111111100000000010000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000000111111110011111111000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000001111111110011111111100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000001111111000101111111100000000000000000000000000000000000000000000000000000000000000000000000010010111010000100001111111000001000100010110001011011111101000000010010000000111111111010000001001111101000101010111011010011110100000010000000000000000000000000000000000000000000000000000000000000000111111110001011001011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110101111111100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001111111110111111110011111111000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011111111111111111110011111111100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011111111111111111110111111111100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011111111111111111110111111111100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001111111110111111110111111111100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010111111110111111111111111111000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000110000101000000001000000011111101100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000101000000001000000000101111110000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111111000000000000000000111111110100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111101000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101000000001000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111100000000001000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111100000000001000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111101000000000000000000111111111100000000000010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111101000000000000100100111111111100000000000100000000000000000100000000000000000000000000000000000000000010000000011000110111010100010110011100010111110010100001001100111110111101001011111111010110011111010000000110001111010111001110110100011000100000000000000000000000000000000000000000000000011000000001000000000000000000000000000010000000010000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111101000000000000000000000000000001111111100000000100000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000001111111101000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111101000000000000000000100000000001111111100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111100000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101000000001000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111111000000000000000000000000000001111111100000000001000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111100000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111111000000000000000000000000000001111111100000000000000000000100000000000000000000000000000000000000000010000000010000111101000000000011100100111111111011111111101111111110100000001001000011110110111100000000000100001111010110011110101000000000001010000000000000000000000000000000000000000000000000000000101111100111110010000000000000000000010111111101100000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000010000011111111101111111111010000000000000000011111111110110000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001111111111111111111000000000000000000010111111110100000000100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000111111111111111111000000000000000000001111111110100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001111111111111111110000000000000000000000111111110100000000100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011111111111111111111000000000000000000010111111110100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011111111111111111111000000000000000000000111111111100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011111111101111111110000000000000000000010111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000011011111110100000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100011110000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111101000000000000000000011111011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111100000000000000000011111111110000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001111111111000000000000000000000111111110100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000001111111110000000000000000000000111111111110000000000000000000000000000000000000000000000000010000000000000000000000000000000000100000000000000000000001111111111000000000000000000010111111110100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001111111111000000000000000000010111111101000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000001111111111100000000000000000010111111101000000000000000000000000000000000000000000000000000010000000010000000000000000000000000100000000000000000000110111111010000000000000000000000111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100111000000110111011111101100000000000000000011100001001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000010010000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000011111011101010111101111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000001111111110111111111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111110111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000001111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111110111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000100011111111110111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000001111111110111111111111111110000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000011011100010000000101000011000100000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;    
    //man greenman8
    parameter [22499:0] greenman8_G3  = 22500'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111011111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111011111111111011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110111111111111111111011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110111111111111111111011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110111111111111111111011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110111111111111111111011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110111111111111111111011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110111111111111111111011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110111111111111111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110111111111111111111011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110011111111101111111011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110111111111000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110111111111000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110111111111000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110111111111000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110111111111000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110111111111000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110111111111000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110111111111000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110111111111000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110111111111000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111101011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter [22499:0] greenman8_G2  = 22500'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111101111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111111100111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111110111111111101111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100011000111111010111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111101111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000111111110111111111011111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111110111111111111101111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111111111111111111111111111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000111111111011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111010111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010011111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111110111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010100000000000010100010011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000011111111101111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111111111111000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111011111111111111111000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111111111111000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111101111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000010000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter [22499:0] greenman8_G1  = 22500'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000001111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010011111111111111111100110000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111001111111110111111101101111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111101111111101111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110111111111110111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111001111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111001111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111001111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111001111111111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010010000000011000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111011111011111111111111111101111101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000111110101111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110111111111001111111001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100111111111011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111110111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111111011111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100110111111101001111110001111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100100000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111101111111110111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111101111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111101111111110111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111101111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111101111111100111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001111111100011110110111111101111111110001111111101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111101111111110111111110111111111100111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111011111111111111111110111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101111111110111111111111111111110111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111101111111111011111111111111111110111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101111111111111111111111111111110111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101111111110011111111011111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101111111111111111111111111111110111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111101111111110011111111101111111100111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101001111110011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110011111111101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100111011100111111110001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111100000000000011111110111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000011111111011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111111000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000111110011001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011101000111111110101011101101111111010001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000001111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000001111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000001111111110111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000001111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000101111111101111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000011111111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111101111111110000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000000000000000000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101111111110000000000000000000000000000001111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111101111111110000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111101111111110000000000000000000000000000000111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111101111111110000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101111111110000000000000000000000000000000111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111101111111110000000000000000000000000000001111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111011111100111111110000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110000000001111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000001111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111110000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111100000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111101111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111101111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111101111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000111111101111111110111111111000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000100000000000000000000000000001110111110111111101011110110100000000000000000000100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    parameter [22499:0] greenman8_G0  = 22500'b000000000000000000000000000000000000000001001111100011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111011111011101101111110011111110001101010100111111100001101110011111111001111111110111011101101011100111111111010111011100111111101010110101100010000000000000000000000000000000000000001111111100011010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000011111111110111111101100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111110011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111110111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000001010000100000000101001111101101111111110011111111001111101010100000000100010011010000000000000100110010110000000001100001001001000000001100000000000000000000000000000000011111111111111111101111111111011111111010000000000000000010000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000111111110111111111100111111101111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111001111111111111111101111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000111111111111111111110011111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000011111111111111111110111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000011111111101111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000111111111111111111110111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101011111111100011111100101111110000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000110100010101011111110010111110000010000000000000000000000000000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000001111111110101111110000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111110111111101000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111110011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111110011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111110011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111111111111110000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000011111111110111111111000000000000000000000000000010000000000000000000100000000000000000000000000000000000000000010000000010000000111010100000110111111010000111111010000001101111111110000010100000000010000000111010010000100011010001001100100110100111000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011111111111111111101100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001111111110101111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011011111111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011111111101111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000000000010011111100111111111100000000000000000010000000000000000000100000000000000000000000000000000000000000010000100010000111101000000010000000001001000111101110000011000000001100110110001111111010001001001000000000100000101001100011100101100101000011111000000000000000000000000000000000000000000000000000001001111100001000010100000000010000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000000000011111111111111111100011111111111111111101000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011111111110111111110111111111111111111111000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010111111111111111111011111110111111111101000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001111111110111111100011111111111111111100010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001111111101111111110011111111111111111100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001111111111111111110111111111011111111111000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011111111111111111110011111111111111111101000000000000000000000000000000000000000000000000000000000000010000000010000000001000000000000000000000000000011111111101111111100111111111111111111101000010000000000000100000000000000000000000000000000000000000010001111010100111101110100110110001010001001111101011100101000000010010000001110000000011111111111000000000111101110001111111100011001101111111001000000000000000000000000000000000000000000000000000000000000000101111000111111110010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110011111111111111111111111111110000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001111111110111111111011111111111111111110000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001111111110111111111111111111111111111110000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000001111111110111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111111111111111111111110000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001111111110011111111101111111110111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111111111111111111010111111111000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001101111100111111101011111000111111010100111010010011111011000000000000000000000000000000000000000000000000000010001000010000000001000000000010000111001111111111111110001000000001000000001110000000011000000001100000000100000000000000000100000000001000000000000010000000000000000000000000000000000000011111110100010111110111111110011111110111111111111101111001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111101111111110111111111111111111111111111110000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111110111111111111111111011111111111111111011111111110000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111110111111111111111110111111111111111111111111111110000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111110111111111111111110011111111111111111111111111110000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111110111111101111111110011111111111111111111111111110000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111110111111111111111101111111110011111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111111111110011111111111111111110111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011000101010000110011111111001111111011111111011000110001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001111011111111111001111011110000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000001111111111111111111111111111101000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000001111111111111111111111111111101000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000001111111111111111111111111111101000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000001111111111111111111111111111101000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000001111111111111111111111111111101000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000001111111111111111111111111111101000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000001111111111111111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111010111111111111011111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000000001111111110011111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000111111110111111111111111111101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110011111111111111111100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000001111111110011111111111111111100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000001111111111011111111111111111101000000000000000000000000000000000000000000000001000000000000010000000000000000000000000000000000000000000000001000000001111111110111111111011111111100000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001111111111111111111111111111110000000000000000000100000000000000000000000000001000000000000010100111010100101101111011000011101100011110101001001111010000000010110000000100000000101000000001011110000101101110001111011100000100101011000000000000000000000000000000000000000000000000000000000000000000001011111000101011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001111111111011111111111111111101000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000111111111001111111111111111101000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000001111111110011111111111111111101000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001111111110011111111111111111101000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000000111111110011111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001111111110111111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111011111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000101110100100111111010001111111010000000000000000000000000000000000000000000000000000000000000010000111011000110001110000000010000000001111111100011011100101011001100000001110000000110000000101100000000110000110000000001100000000101000001001000010000000000000000000000000000000000000000000000000101111010000000000011111110101111111110000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000000000011111111100000000000011111111111111111101000000001000000000100000000000000000000000000001000000000000010000000000000000000000000000000000000000000000011111111001000000000111111111011111111101000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011111111110000000000111111111111111111101000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001111111100000000000111111111111111111101000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011111111110000000000111111111111111111001000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001111111111000000100111111111111111111101000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000011011111110100000000111111111111111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100101001111100110110001001111111111110111110001000000000000000000000000000000000000000000000000000010000000011000110111000010000110011010000000011000011101010111110011011011101000000000111011111111000010100110001010001001001100110100111000100000000000000000000000000000000000000000000000000000000000000000001111111111000000000101110111110111111001000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001111111111000000000101111111111111111111100000000100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000001111111110100000000101111111111111111110000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000001111111111100000000101111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111100000000101111111011111111110000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000000111111111000000000101111111111111111110000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000001111111111100000000101111111111111111101000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000000000000000000001111111110100000000001111111100111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001111100010001101111101011100000000111001000011000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000110110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111101010111110111111100000000000000000000000000000001111111010100000000000000000000000000000000000000000010000000010000000000000000000000000000011111111110111111101111111110000000000000000000000000000000111111110010000000000000000000000000000000000000000010000000000000000000000000000000000000011111111110111111111111111111100000000000000000000000000000111111111000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111111111111110111111111000000000000000000000000000001111111110000000000000000000000000000000000000000000010000000000000000000000000000000000000011111111111111111111111111111100000000000000000010000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110111111110111111111100000000000000000000000000001111111110000000000000000000000000000000000000000000010000000000000000000000000000000000000001111111110111111111111111111100000000000000000000000000001111111111100000000000000000000000000000000000000000010000000010000000000000000000000000000001111111110011111111111111111100000000000000000010000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011100000001010001011100001000110000000011111111010000000001111101111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000010000000001010000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000111111111110000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000101111111100000000001111111111000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000000000000000000000000101111111100000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111100000000001111111111000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000000000000000000000000101111111100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000001111111111000000001111111111100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000001000000001000000000000000000101111111101000000000011111110010000000000000000000000000001000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000001111111010111111101101111110110000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000010000010000010000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011111111111111101101111111110000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111110000000000000000000000000000000010000000000000000000000000000000000000000000000001000000000000000000000000000000000000010111111111111111111111111111010000000000000000000000000000000010000000000000000001000000000000000000000000000001000000000000000000000000000000000000001111111111111111111111111111110000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111110000000100000000000000000000000010000000000000000000000000000000000000000000000001000000000000000000000000000000000000001111111110111111111011111111110000000000000000000000000001000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000001111111111111111111011111111110000000000000000000000000000000010000000010000000000000000000000000000000000000000000000000000000000000000000100000000011111111111111111111111111111110000000000000000000000000000000011111110001000011101111110010111101111011111111011111111000111111110110110101101111111000110111100001111101001110110001111111101100100000111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;    

    //-----640*480---------------------------------
    parameter H_ACTIVE = 640;
    parameter H_SYNC = 96;
    parameter H_BP = 48;
    parameter H_FP = 16;
    parameter H_WHOLE = 800;
    parameter V_ACTIVE = 480;
    parameter V_SYNC = 2;
    parameter V_BP = 33;
    parameter V_FP = 10;
    parameter V_WHOLE = 525;
  
    reg  [30:0] counter, next_counter;
    reg  [9:0]  counth, countv, px, py;
    wire [9:0]  next_counth, next_countv;
    reg  [3:0]  next_vgaRed, next_vgaBlue, next_vgaGreen;
    reg  [20:0] tmp;
    
    assign Hsync = (counth < H_SYNC)?1'b1:1'b0;
    assign Vsync = (countv < V_SYNC)?1'b1:1'b0;
    assign next_counth = (counth == H_WHOLE-1)?11'd0:counth+1;
    assign next_countv = (counth == H_WHOLE-1)?((countv==V_WHOLE-1)?11'd0:countv+1):countv;
    
    always@(*) begin
        if(counth >= (H_SYNC+H_BP) && counth < (H_SYNC+H_BP+H_ACTIVE) && countv >= (V_SYNC+V_BP) && countv < (V_SYNC+V_BP+V_ACTIVE)) begin
            px = counth-(H_SYNC+H_BP);
            py = countv-(V_SYNC+V_BP);
            
            //----------------The car traffic light part---------------------
            if(px >= 50 && px <150 && py>=50 && py<150) begin  //Red light(light[2])
                tmp = 9999-((py-50)*100+px-50);
                if(car_R==0) begin  //black light
                    next_vgaRed     = 4'b0000; 
                    next_vgaBlue    = 4'b0000;
                    next_vgaGreen[3]   = black_G3[tmp];
                    next_vgaGreen[2:0] = 3'b000;
                end
                else begin //red light on
                    next_vgaRed[3]     = red_R3[tmp]; 
                    next_vgaRed[2:0]   = {{3{next_vgaRed[3]}}};
                    next_vgaGreen[3]   = red_G3[tmp];
                    next_vgaBlue    = 4'b0000;
                    next_vgaGreen[2:0] = 3'b000;
                end
            end
            else if(px >= 150 && px <250 && py>=50 && py<150) begin  //Yellow light (light[1])
                tmp = 9999-((py-50)*100+px-150);
                if(car_Y==0) begin  //black light
                    next_vgaRed     = 4'b0000; 
                    next_vgaBlue    = 4'b0000;
                    next_vgaGreen[3]   = black_G3[tmp];
                    next_vgaGreen[2:0] = 3'b000;
                end
                else begin //yellow light on
                    next_vgaBlue       = 4'b0000;
                    next_vgaGreen[3]   = 1'b1;
                    next_vgaGreen[2]   = green_G2[tmp];
                    next_vgaGreen[1:0] = {{2{next_vgaGreen[2]}}};
                    next_vgaRed        = {{4{next_vgaGreen[2]}}};
                end            
            end
            else if(px >= 250 && px <350 && py>=50 && py<150) begin  //Green light  (light[0])
                tmp = 9999-((py-50)*100+px-250);
                if(car_G==0) begin  //black light
                    next_vgaRed     = 4'b0000; 
                    next_vgaBlue    = 4'b0000;
                    next_vgaGreen[3]   = black_G3[tmp];
                    next_vgaGreen[2:0] = 3'b000;
                end
                else begin //green light on
                    next_vgaBlue       = 4'b0000;
                    next_vgaRed        = 4'b0000;
                    next_vgaGreen[3]   = 1'b1;
                    next_vgaGreen[2]   = green_G2[tmp];
                    next_vgaGreen[1:0] = {{2{next_vgaGreen[2]}}};
                end                
            end
            //----------------The man traffic light part---------------------
            else if(px >= 450 && px <600 && py>=50 && py<200) begin  //Red man
                tmp = 22499-((py-50)*150+px-450);
                if(man_R==0) begin  //red man light off -> black
                    next_vgaBlue       = 4'b0000;
                    next_vgaRed        = 4'b0000;
                    next_vgaGreen      = 4'b0000;
                end
                else begin //red man light on
                    next_vgaBlue       = 4'b0000;
                    next_vgaGreen      = 4'b0000;
                    next_vgaRed[3]     = redman_R3[tmp];
                    next_vgaRed[2]     = redman_R2[tmp];
                    next_vgaRed[1]     = redman_R1[tmp];
                    next_vgaRed[0]     = redman_R0[tmp];
                end                
            end            
            else if(px >= 450 && px <600 && py>=200 && py<350) begin  //Green man
                tmp = 22499-((py-200)*150+px-450);
                if(man_G_ID==1) begin  //green man 1
                    next_vgaBlue       = 4'b0000;
                    next_vgaRed        = 4'b0000;
                    next_vgaGreen[3]   = greenman1_G3[tmp];
                    next_vgaGreen[2]   = greenman1_G2[tmp];
                    next_vgaGreen[1]   = greenman1_G1[tmp];
                    next_vgaGreen[0]   = greenman1_G0[tmp];                    
                end
                else if(man_G_ID==2) begin  //green man 1
                    next_vgaBlue       = 4'b0000;
                    next_vgaRed        = 4'b0000;
                    next_vgaGreen[3]   = greenman2_G3[tmp];
                    next_vgaGreen[2]   = greenman2_G2[tmp];
                    next_vgaGreen[1]   = greenman2_G1[tmp];
                    next_vgaGreen[0]   = greenman2_G0[tmp];                    
                end
                else if(man_G_ID==3) begin  //green man 1
                    next_vgaBlue       = 4'b0000;
                    next_vgaRed        = 4'b0000;
                    next_vgaGreen[3]   = greenman3_G3[tmp];
                    next_vgaGreen[2]   = greenman3_G2[tmp];
                    next_vgaGreen[1]   = greenman3_G1[tmp];
                    next_vgaGreen[0]   = greenman3_G0[tmp];                    
                end
                else if(man_G_ID==4) begin  //green man 1
                    next_vgaBlue       = 4'b0000;
                    next_vgaRed        = 4'b0000;
                    next_vgaGreen[3]   = greenman4_G3[tmp];
                    next_vgaGreen[2]   = greenman4_G2[tmp];
                    next_vgaGreen[1]   = greenman4_G1[tmp];
                    next_vgaGreen[0]   = greenman4_G0[tmp];                    
                end
                else if(man_G_ID==5) begin  //green man 1
                    next_vgaBlue       = 4'b0000;
                    next_vgaRed        = 4'b0000;
                    next_vgaGreen[3]   = greenman5_G3[tmp];
                    next_vgaGreen[2]   = greenman5_G2[tmp];
                    next_vgaGreen[1]   = greenman5_G1[tmp];
                    next_vgaGreen[0]   = greenman5_G0[tmp];                    
                end
                else if(man_G_ID==6) begin  //green man 1
                    next_vgaBlue       = 4'b0000;
                    next_vgaRed        = 4'b0000;
                    next_vgaGreen[3]   = greenman6_G3[tmp];
                    next_vgaGreen[2]   = greenman6_G2[tmp];
                    next_vgaGreen[1]   = greenman6_G1[tmp];
                    next_vgaGreen[0]   = greenman6_G0[tmp];                    
                end
                else if(man_G_ID==7) begin  //green man 1
                    next_vgaBlue       = 4'b0000;
                    next_vgaRed        = 4'b0000;
                    next_vgaGreen[3]   = greenman7_G3[tmp];
                    next_vgaGreen[2]   = greenman7_G2[tmp];
                    next_vgaGreen[1]   = greenman7_G1[tmp];
                    next_vgaGreen[0]   = greenman7_G0[tmp];                    
                end
                else if(man_G_ID==8) begin  //green man 1
                    next_vgaBlue       = 4'b0000;
                    next_vgaRed        = 4'b0000;
                    next_vgaGreen[3]   = greenman8_G3[tmp];
                    next_vgaGreen[2]   = greenman8_G2[tmp];
                    next_vgaGreen[1]   = greenman8_G1[tmp];
                    next_vgaGreen[0]   = greenman8_G0[tmp];                    
                end
                else begin //green man light off
                    next_vgaBlue       = 4'b0000;
                    next_vgaRed        = 4'b0000;
                    next_vgaGreen      = 4'b0000;
                end                
            end               
            else begin
                tmp = 0;
                next_vgaRed     = 4'b1111;
                next_vgaGreen   = 4'b1111;
                next_vgaBlue    = 4'b1111;                 
            end
        end
        
        else begin
            tmp = 0;
            next_vgaRed = 4'b0000;
            next_vgaGreen = 4'b0000;
            next_vgaBlue = 4'b0000; 
        end
    end
    
    
    always@(posedge clk or posedge rst) begin
        if(rst) begin
            counter <= 0;
            vgaRed  <= 4'b0;
            vgaGreen<= 4'b0;
            vgaBlue <= 4'b0;
            counth  <= 0;
            countv  <= 0;
        end
        else begin
            counter <= next_counter;
            vgaRed  <= next_vgaRed  ;
            vgaGreen<= next_vgaGreen;
            vgaBlue <= next_vgaBlue ;
            counth  <= next_counth ;
            countv  <= next_countv;
        end
    end
    
endmodule
